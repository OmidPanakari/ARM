module InstructionMemory (
    address,
    instruction
);
    input [31:0] address;
    output [31:0] instruction;
    reg [31:0] mem [0:1023];
    integer i;

    initial begin
        for (i = 0; i < 1024; i = i + 1) begin
            mem[i] = 32'd0;
        end
        mem[0] = 32'b1110_00_1_1101_0_0000_0000_000000010100; // MOV    R0,#20  =>  R0=20
        mem[1] = 32'b1110_00_1_1101_0_0000_0001_101000000001; // MOV    R1,#4096    =>  R1=4096
        mem[2] = 32'b1110_00_1_1101_0_0000_0010_000100000011; // MOV    R2,#0xC0000000  =>  R2=-1073741824
        mem[3] = 32'b1110_00_0_0100_1_0010_0011_000000000010; // ADDS   R3,R2,R2    =>  R3=-2147483648
        mem[4] = 32'b1110_00_0_0101_0_0000_0100_000000000000; // ADC    R4,R0,R0    =>  R4=41
        mem[5] = 32'b1110_00_0_0010_0_0100_0101_000100000100; // SUB    R5,R4,R4,LSL #2 => R5=-123
        mem[6] = 32'b1110_00_0_0110_0_0000_0110_000010100000; // SBC    R6,R0,R0,LSR #1 => R6=10
        mem[7] = 32'b1110_00_0_1100_0_0101_0111_000101000010; // ORR    R7,R5,R2,ASR #2 => R7=-123
        mem[8] = 32'b1110_00_0_0000_0_0111_1000_000000000011; // AND    R8,R7,R3    =>  R8=-2147483648
        mem[9] = 32'b1110_00_0_1111_0_0000_1001_000000000110; // MVN    R9,R6   =>  R9=-11
        mem[10] = 32'b1110_00_0_0001_0_0100_1010_000000000101; // EOR   R10,R4,R5   =>  R10=-84
        mem[11] = 32'b1110_00_0_1010_1_1000_0000_000000000110; // CMP   R8,R6
        mem[12] = 32'b0001_00_0_0100_0_0001_0001_000000000001; // ADDNE R1,R1,R1    =>  R1=8192
        mem[13] = 32'b1110_00_0_1000_1_1001_0000_000000001000; // TST   R9,R8
        mem[14] = 32'b0000_00_0_0100_0_0010_0010_000000000010; // ADDEQ R2,R2,R2    =>  R2=-1073741824
        mem[15] = 32'b1110_00_1_1101_0_0000_0000_101100000001; // MOV   R0,#1024    =>  R0=1024
        mem[16] = 32'b1110_01_0_0100_0_0000_0001_000000000000; // STR   R1,[R0],#0  =>  Mem[1024]=8192
        mem[17] = 32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR    R11,[R0],#0 =>  R11=8192
        mem[18] = 32'b1110_01_0_0100_0_0000_0010_000000000100; //STR	
        mem[19] = 32'b1110_01_0_0100_0_0000_0011_000000001000; //STR
        mem[20] = 32'b1110_01_0_0100_0_0000_0100_000000001101; //STR
        mem[21] = 32'b1110_01_0_0100_0_0000_0101_000000010000; //STR
        mem[22] = 32'b1110_01_0_0100_0_0000_0110_000000010100; //STR	
        mem[23] = 32'b1110_01_0_0100_1_0000_1010_000000000100; //LDR
        mem[24] = 32'b1110_01_0_0100_0_0000_0111_000000011000; //STR
        mem[25] = 32'b1110_00_1_1101_0_0000_0001_000000000100; //MOV
        mem[26] = 32'b1110_00_1_1101_0_0000_0010_000000000000; //MOV
        mem[27] = 32'b1110_00_1_1101_0_0000_0011_000000000000; //MOV
        mem[28] = 32'b1110_00_0_0100_0_0000_0100_000100000011; //ADD
        mem[29] = 32'b1110_01_0_0100_1_0100_0101_000000000000; //LDR
        mem[30] = 32'b1110_01_0_0100_1_0100_0110_000000000100; //LDR
        mem[31] = 32'b1110_00_0_1010_1_0101_0000_000000000110; //CMP
        mem[32] = 32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGT
        mem[33] = 32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGT
        mem[34] = 32'b1110_00_1_0100_0_0011_0011_000000000001; //ADD
        mem[35] = 32'b1110_00_1_1010_1_0011_0000_000000000011; //CMP
        mem[36] = 32'b1011_10_1_0_111111111111111111110111   ; //BLT
        mem[37] = 32'b1110_00_1_0100_0_0010_0010_000000000001; //ADD
        mem[38] = 32'b1110_00_0_1010_1_0010_0000_000000000001; //CMP	
        mem[39] = 32'b1011_10_1_0_111111111111111111110011   ; //BLT
        mem[40] = 32'b1110_01_0_0100_1_0000_0001_000000000000; //LDR
        mem[41] = 32'b1110_01_0_0100_1_0000_0010_000000000100; //LDR
        mem[42] = 32'b1110_01_0_0100_1_0000_0011_000000001000; //LDR
        mem[43] = 32'b1110_01_0_0100_1_0000_0100_000000001100; //LDR
        mem[44] = 32'b1110_01_0_0100_1_0000_0101_000000010000; //LDR
        mem[45] = 32'b1110_01_0_0100_1_0000_0110_000000010100; //LDR
        mem[46] = 32'b1110_10_1_0_111111111111111111111111   ; //B	

    end
    
    assign instruction = mem[(address >> 2)];
endmodule