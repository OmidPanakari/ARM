module Execution (
    clk,
    rst,
    pc
);
    input clk, rst;
    input [31:0] pc;
endmodule